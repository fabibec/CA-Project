----------------------------------------------------------------------------------
-- Engineers: Fabian Becker, Nicolas Koch
-- 
-- Create Date: 05/22/2025 03:08:36 PM
-- Design Name: 
-- Module Name: as_core - arch
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity as_core is
    generic (
        UART_BAUDRATE_DIVISOR: integer := 651;
        UART_NUM_DATA_BITS: integer := 8;
        CONTROL_MS_DIVISOR: integer := 100_000;
        CONTROL_POWER_UP_TIME : integer := 250; -- 250 ms power-up delay
        CONTROL_FIRST_READING_TIME : integer := 100; -- 100 ms first reading delay
        -- the sensor checks if tx is high every 49 ms and then proceeds to measrue or not
        -- so worst case time can be 2x interval!!
        CONTROL_CALIBRATION_TIME : integer := 49; -- 49 ms calibration cycle
        CONTROL_RANGE_READING_TIME : integer := 49 -- 49 ms range reading time
    );
    port ( 
        -- AXI 
        i_clk: in std_logic;
        i_reset: in std_logic;
        
        -- GCSR
        i_ap_start: in std_logic;
        o_ap_idle: out std_logic; -- async, register when ad_done -> 1, on i_ap_start or reset or restart = 0 
        o_ap_done: out std_logic; -- ad_done    
        i_auto_restart: in std_logic; 
        
        -- SCSR0
        o_powerup_done: out std_logic;
        o_calib_done: out std_logic;
        o_read_valid: out std_logic; -- no ad_error, uart can be ignored, updated/set on done
        i_reset_ip: in std_logic; 
        i_freeze_ip: in std_logic; -- # TODO ONLY accept freeze if no reset in progess!!!
 
        -- DIST0
        o_dist_in: out std_logic_vector(7 downto 0); -- ad_data, updated/set on done
        o_dist_char_1: out std_logic_vector(7 downto 0); -- ad_char 1
        o_dist_char_2: out std_logic_vector(7 downto 0); -- ad_char 2 
        o_dist_char_3: out std_logic_vector(7 downto 0);
 
       -- UCSR Signals
       o_ur_error: out std_logic; -- ur_error, updated async, 1 if at least on error occured during current measurement reading, cleared on start 
       o_ur_data: out std_logic_vector(7 downto 0); -- ur_data, updated async, cleared on start
 
       -- ADSR Signals
       o_ad_error: out std_logic; -- ad_error, updated/set on done
       o_ad_err_pos: out std_logic_vector(5 downto 0); -- ad_err_pos, updated/set on done
       o_ad_err_char: out std_logic_vector(7 downto 0); -- ad_err_char, updated/set on done
       
       -- I/Os
       i_rx: in std_logic;
       o_tx: out std_logic
    );
end as_core;

architecture arch of as_core is

    -- Control Timer 
    component control_timer is
    generic (
        MS_DIVISOR : integer := 100_000; -- 1 ms @ 100 MHz
        POWER_UP_TIME : integer := 250; -- 250 ms power-up delay
        FIRST_READING_TIME : integer := 100; -- 100 ms first reading delay
        CALIBRATION_TIME : integer := 49; -- 49 ms calibration cycle
        RANGE_READING_TIME : integer := 49 -- 49 ms range reading time
    );
    port (
        i_clk : in std_logic;
        i_reset : in std_logic;
        i_enable: in std_logic; 
        i_reset_timer: in std_logic;
        o_done : out std_logic := '0';
        o_powerup_done : out std_logic := '0';
        o_config_done : out std_logic := '0';
        o_init_done : out std_logic := '0'
        
    );
    end component;

    -- Counter for Baudrate generation
    component baud_rate_generator is
        generic (
            DIVISOR : integer
        );
        port (
            i_enable: in std_logic;
            i_clk: in std_logic;  
            i_reset: in std_logic;
            o_tick: out std_logic
        );
    end component;
    
    -- UART Receiver for sensor data
    component uart_receiver is
        generic (
            OVERSAMPLING_TICK_START: integer;
            OVERSAMPLING_TICK_DATA: integer;
            N_DATA_BITS: integer
        );
        port(
            -- I/Os 
            i_rx: in std_logic; -- UART Receive
            
            -- UART Receiver control
            i_enable: in std_logic; 
            i_tick: in std_logic; -- generated by the baud rate generator
            i_clk: in std_logic;
            i_reset: in std_logic;
            
            -- Baud rate control
            o_baud_enable: out std_logic; -- enable baud rate generator
            
            -- Output
            o_done: out std_logic;
            o_data: out unsigned(7 downto 0);
            o_error: out std_logic;
            
            -- Debug 
            o_sample: out std_logic
        );
    end component;
    
    -- ASCII Decoder to convert UART data to 1 byte number
    component ascii_decoder is
        port(
            -- Input
            i_enable: in std_logic;
            i_uart_char: in unsigned(7 downto 0);
            i_uart_char_ready: in std_logic;
            i_sensor_cycle_done: in std_logic;
            i_clk: in std_logic;
            i_reset: in std_logic;
            
            -- Output
            o_start: out std_logic;
            o_done: out std_logic;
            o_data: out unsigned(7 downto 0);
            o_error: out std_logic;
            o_error_pos: out std_logic_vector(5 downto 0);
            o_error_char: out std_logic_vector(7 downto 0);
            
            -- Debug
            o_digit: out std_logic_vector(7 downto 0);
            o_digit_ready: out std_logic;
            o_chars: out std_logic_vector(3 downto 0)
        );
    end component;
    
    signal ap_start_stage1, ap_start_stage2: std_logic := '0';
    signal global_enable: std_logic;
    
    signal global_reset: std_logic := '0';
    
    signal sensor_enable: std_logic;
    
    signal ctl_reset_timer: std_logic;
    signal ctl_enable: std_logic;
    signal ctl_done: std_logic;
    signal ctl_powerup_done: std_logic;
    signal ctl_calib_done: std_logic;
    
    signal bd_gen_enable: std_logic;
    signal bd_gen_tick: std_logic;
    
    signal ur_baud_enable: std_logic;
    signal ur_done: std_logic;
    signal ur_data: unsigned(7 downto 0);
    signal ur_error: std_logic;
    
    signal ad_start: std_logic;
    signal ad_done: std_logic;
    signal ad_data: unsigned(7 downto 0);
    signal ad_error, ad_error_reg: std_logic;
    signal ad_err_pos, ad_err_pos_reg: std_logic_vector(5 downto 0);
    signal ad_err_char, ad_err_char_reg: std_logic_vector(7 downto 0);
    signal ad_digit_ready: std_logic;
    signal ad_digit: std_logic_vector(7 downto 0);
    
    signal ad_dist_in_reg: std_logic_vector(7 downto 0) := (others => '0');
    signal ad_dist_char_1_reg: std_logic_vector(7 downto 0) := (others => '0');
    signal ad_dist_char_2_reg: std_logic_vector(7 downto 0) := (others => '0');
    signal ad_dist_char_3_reg: std_logic_vector(7 downto 0) := (others => '0');
    signal ad_digit_index: unsigned(1 downto 0) := (others => '0'); -- (0-3)
    
    signal read_valid_reg: std_logic := '0';
    signal update_window: std_logic := '0';
    
    -- Debug
    signal ur_sample: std_logic;
    signal ad_chars: std_logic_vector(3 downto 0);

begin
    -- Write big ass testbench
    
    CONTROL_TIMER_INST: control_timer
        generic map (
            MS_DIVISOR => CONTROL_MS_DIVISOR,
            POWER_UP_TIME => CONTROL_POWER_UP_TIME,
            FIRST_READING_TIME => CONTROL_FIRST_READING_TIME,
            CALIBRATION_TIME => CONTROL_CALIBRATION_TIME,
            RANGE_READING_TIME => CONTROL_RANGE_READING_TIME
        )
        port map (
            i_clk => i_clk,
            i_reset => global_reset,
            i_enable => ctl_enable,
            i_reset_timer => ctl_reset_timer,
            o_done => ctl_done,
            o_powerup_done => ctl_powerup_done,
            o_config_done => ctl_calib_done,
            o_init_done => open
        );

    -- Instantion of Baudrate Generator
    BAUD_GEN_INST: baud_rate_generator
        generic map (
            DIVISOR => UART_BAUDRATE_DIVISOR
        )
        port map (
            i_enable => bd_gen_enable,
            i_clk => i_clk,
            i_reset => global_reset,
            o_tick => bd_gen_tick
        );
        
    -- Instantion of UART Receiver
    UART_RECEIVER_INST: uart_receiver
        generic map (
            OVERSAMPLING_TICK_START => 7,
            OVERSAMPLING_TICK_DATA => 15,
            N_DATA_BITS => UART_NUM_DATA_BITS
        )
        port map (
            -- I/Os 
            i_rx => i_rx,
            
            -- UART Receiver control
            i_enable => sensor_enable,
            i_tick => bd_gen_tick,
            i_clk => i_clk,
            i_reset => global_reset,
            
            -- Baud rate control
            o_baud_enable => ur_baud_enable,
            
            -- Output
            o_done => ur_done,
            o_data => ur_data,
            o_error => ur_error,
            
            -- Debug 
            o_sample => ur_sample
        );
    
    -- Instantion of ASCII Decoder
    ASCII_DECODER_INST: ascii_decoder
        port map (
            -- Input
            i_enable => sensor_enable,
            i_uart_char => ur_data,
            i_uart_char_ready => ur_done,
            i_sensor_cycle_done => ctl_done,
            i_clk => i_clk,
            i_reset => global_reset,
            
            -- Output
            o_start => ad_start,
            o_done => ad_done,
            o_data => ad_data,
            o_error => ad_error,
            o_error_pos => ad_err_pos,
            o_error_char => ad_err_char,
            
            -- Debug
            o_digit => ad_digit,
            o_digit_ready => ad_digit_ready,
            o_chars => ad_chars
        );

    -- ad_done will be stretched interally to one more clock cycle unless the ip is frozen
    -- the strected output will serve as an enable signal to make sure the synchronous resets are excuted properly after ap_done is high
    AP_START_STRETCH_PROC: process(i_clk)
    begin
        if (i_clk'event and i_clk = '1') then
            if global_reset = '1' then
                ap_start_stage1 <= '0';
                ap_start_stage2 <= '0';
            elsif i_freeze_ip = '0' then
                ap_start_stage1 <= i_ap_start;
                ap_start_stage2 <= ap_start_stage1;
            end if;
        end if;
    end process;
    
    -- Concurrent signal assignments
    global_reset <= i_reset or i_reset_ip;
    global_enable <= ap_start_stage1 or ap_start_stage2;
    
    ctl_enable <= not i_freeze_ip and global_enable; -- stretch ap_start by 1 clock cycle in order to enable timer reset
    ctl_reset_timer <= ad_done; 
    
    sensor_enable <= ctl_enable and ctl_calib_done;
    
    bd_gen_enable <= sensor_enable and ur_baud_enable;

    -- Output assignments
    o_ap_idle <= not i_ap_start;
    
    o_powerup_done <= ctl_powerup_done;
    o_calib_done <= ctl_calib_done;
    o_ap_done <= ad_done;

    -- one clock of stable output during the done signal it not enough for software to read the results
    -- therefor this process will keep the distance and ascii decoder outputs stable, updating this data is only allowed
    -- after the ascii decoder starts and until the done signal ends. So even if there is a timeout error the system is able to update for one clock
    OUTPUT_UPDATE_PROC: process (i_clk)
    begin 
        if (i_clk'event and i_clk = '1') then
            if global_reset = '1' or ad_start = '1' then
                read_valid_reg <= '0';
                update_window <= '0';
                
                ad_dist_in_reg <= (others => '0');
                ad_dist_char_1_reg <= (others => '0');
                ad_dist_char_2_reg <= (others => '0');
                ad_dist_char_3_reg <= (others => '0');
                ad_digit_index <= (others => '0');
                
                ad_error_reg <= '0';
                ad_err_pos_reg <= (others => '0');
                ad_err_char_reg <= (others => '0');
                
                if ad_start = '1' then 
                   update_window <= '1';
                end if;
            elsif i_freeze_ip = '0' then                
                if update_window = '1' then
                    -- Distance in inches
                    ad_dist_in_reg <= std_logic_vector(ad_data);
                    -- Distance Chars 
                    if ad_digit_ready = '1' then
                        case ad_digit_index is
                            when "00" =>
                                ad_dist_char_1_reg <= ad_digit;
                            when "01" =>
                                ad_dist_char_2_reg <= ad_digit;
                            when "10" =>
                                ad_dist_char_3_reg <= ad_digit;
                            when others =>
                                null;
                        end case;
    
                        if ad_digit_index < 2 then
                            ad_digit_index <= ad_digit_index + 1;
                        end if;
                    end if;
                    -- ASCII Decoder
                    ad_error_reg <= ad_error;
                    ad_err_pos_reg <= ad_err_pos;
                    ad_err_char_reg <= ad_err_char;    
                    -- Read is valid after done
                    if ad_done = '1' then
                        read_valid_reg <= '1';
                    end if;
                    -- Close update window
                    if ad_done = '1' then
                        update_window <= '0';
                    end if;
                end if;         
            end if;
        end if;
    end process;
    
    o_read_valid <= read_valid_reg;
    
    o_dist_in <= ad_dist_in_reg;
    o_dist_char_1 <= ad_dist_char_1_reg;
    o_dist_char_2 <= ad_dist_char_2_reg;
    o_dist_char_3 <= ad_dist_char_3_reg;
    
    o_ad_error <= ad_error_reg;
    o_ad_err_char <= ad_err_char_reg;
    o_ad_err_pos <= ad_err_pos_reg;
    
    o_ur_data <= std_logic_vector(ur_data);
    o_ur_error <= ur_error;
    
    o_tx <= i_ap_start or i_auto_restart;

end arch;
