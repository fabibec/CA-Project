----------------------------------------------------------------------------------
-- Engineer: Fabian Becker, Nicolas Koch
-- 
-- Create Date: 05/09/2025 08:01:52 PM
-- Design Name: 
-- Module Name: uart_receiver - arch
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity uart_receiver is
    generic (
        OVERSAMPLING_TICK_START : integer := 7;
        OVERSAMPLING_TICK_DATA  : integer := 15;
        N_DATA_BITS             : integer := 8
    );
    port(
        -- I/Os 
        i_rx: in std_logic; -- UART Receive
        
        -- UART Receiver control
        i_enable: in std_logic; 
        i_tick: in std_logic; -- generated by the baud rate generator
        i_clk: in std_logic;
        i_reset: in std_logic;
        
        -- Baud rate control
        o_baud_enable: out std_logic; -- enable baud rate generator
        
        -- Output
        o_done: out std_logic;
        o_data: out unsigned((N_DATA_BITS - 1) downto 0);
        o_error: out std_logic;
        
        -- Debug 
        o_sample: out std_logic
    );
end uart_receiver;

architecture arch of uart_receiver is
    type state_type is (idle, start, data, stop); 
    
    signal state, next_state: state_type; 
    signal ticks_reg, ticks_next: unsigned (3 downto 0) := (others => '0'); -- ticks
    signal baud_enable_reg, baud_enable_next : std_logic := '0';
    signal bits_reg, bits_next: unsigned (3 downto 0) := (others => '0'); -- # data bits
    signal data_reg, data_next: unsigned ((N_DATA_BITS - 1) downto 0) := (others => '0'); -- uart rx register
    
    signal error_next: std_logic := '0';
    signal done_next: std_logic := '0';
    
begin

    NSTATEPROC: process(
        state, i_rx, i_tick, i_enable, ticks_reg, bits_reg, data_reg, baud_enable_reg
    )
    begin
        -- Default values
        next_state <= state;
        ticks_next <= ticks_reg;
        bits_next <= bits_reg;
        data_next <= data_reg;
        baud_enable_next <= baud_enable_reg;
        done_next <= '0';
        error_next <= '0';
        o_sample <= '0';
            
        if i_enable = '1' then
            case state is
                when idle =>
                    if (i_rx'event and i_rx = '0' and i_enable = '1') then
                        next_state <= start;
                        ticks_next <= (others => '0');
                        data_next <= (others => '0');
                        baud_enable_next <= '1';  -- start baud
                    end if;
    
                when start =>
                    if i_tick = '1' then 
                        if ticks_reg = OVERSAMPLING_TICK_START then
                            next_state <= data;
                            ticks_next <= (others => '0');
                            bits_next <= (others => '0');
                            o_sample <= '1';
                        else
                            ticks_next <= ticks_reg + 1;
                        end if;
                    end if;
    
                when data =>
                    if i_tick = '1' then 
                        if ticks_reg = OVERSAMPLING_TICK_DATA then
                            ticks_next <= (others => '0');
                            o_sample <= '1';
                            data_next <= i_rx & data_reg(7 downto 1); -- LSB first
                            --data_next <= data_reg(6 downto 0) & i_rx; -- MSB first
    
                            if bits_reg = (N_DATA_BITS - 1) then
                                next_state <= stop;
                            else
                                bits_next <= bits_reg + 1;
                            end if;
                        else 
                            ticks_next <= ticks_reg + 1;
                        end if;
                    end if;
    
                when stop =>
                    if i_tick = '1' then 
                        if ticks_reg = OVERSAMPLING_TICK_DATA then
                            o_sample <= '1';
                            if (i_rx /= '1') then
                                error_next <= '1';
                            end if;
                            next_state <= idle;
                            done_next <= '1';
                            baud_enable_next <= '0';
                        else
                            ticks_next <= ticks_reg + 1;
                        end if;
                    end if;
    
                when others =>
                    null;
            end case;
        end if;
    end process;

    
    STATEPROC: process(i_clk)
    begin
        if (i_clk'event and i_clk = '1') then
            if i_reset = '1' then
                state <= idle;
                ticks_reg <= (others => '0');
                bits_reg <= (others => '0');
                data_reg <= (others => '0');
                baud_enable_reg <= '0';
                o_error <= '0';
                o_done <= '0';
            else
                if i_enable = '1' then
                    state <= next_state;
                    ticks_reg <= ticks_next;
                    bits_reg <= bits_next;
                    data_reg <= data_next;
                    baud_enable_reg <= baud_enable_next;
                    o_done <= done_next;
                    o_error <= error_next;
                end if;
            end if;
        end if;
    end process;
    
    o_data <= data_reg;
    o_baud_enable <= baud_enable_reg;

end arch;